module driver (
	output wire r, g, b
);

	assign {r, g, b} = 3'b111;

endmodule
