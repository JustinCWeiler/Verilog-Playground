module SB_HFOSC #(
	parameter CLKHF_DIV = "0b00"
)
(
	input logic CLKHFEN, CLKHFPU,
	output logic CLKHF
);
endmodule
