module driver (
	output logic r, g, b
);

	assign {r, g, b} = 3'b111;

endmodule
